module scoreDisplay(input logic clk, reset,
								input logic [8:0] score,
								output logic leftDigitTransBase, rightDigitTransBase,
								output logic [6:0] seg,
								output logic );
	
	//Alternate LEDs at clk/(32768)=1220 Hz
	logic [16:0] counter; //16-bit counter
	logic switch; //LED group to drive (0 or 1)
	assign switch = counter[16]; //highest bit of counter
	always_ff @(posedge clk)
		counter <= counter + 1;
	//Only one transistor base low at a time
	assign leftDigitTransBase = switch;
	assign rightDigitTransBase = ~switch;
	//Switch to 7-segment display decoder
	logic [3:0] leftDigit;
	assign leftDigit = score/10;
	logic [3:0] rightDigit;
	assign rightDigit = score%10;
	hexto7seg dispDecoder(clk,,seg);
endmodule

//Module that decodes hexadecimal value to 7- segment display
module hexto7seg(input logic clk, input logic [3:0] hex, output logic [6:0] seg);
	//Common logic-high anode, output is cathode value
	//Logic-low output indicates turning segment
	always_comb begin
		case (hex)
			4'h0: seg <= 7'b1000000;
			4'h1: seg <= 7'b1111001;
			4'h2: seg <= 7'b0100100;
			4'h3: seg <= 7'b0110000;
			4'h4: seg <= 7'b0011001;
			4'h5: seg <= 7'b0010010;
			4'h6: seg <= 7'b0000010;
			4'h7: seg <= 7'b1111000;
			4'h8: seg <= 7'b0000000;
			4'h9: seg <= 7'b0011000;
			4'hA: seg <= 7'b0001000; //A
			4'hB: seg <= 7'b0000011; //b
			4'hC: seg <= 7'b1000110; //C
			4'hD: seg <= 7'b0100001; //d
			4'hE: seg <= 7'b0000110; //E
			4'hF: seg <= 7'b0001110; //F
		endcase
	end
endmodule
